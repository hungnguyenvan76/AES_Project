`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/01/2025 08:43:40 PM
// Design Name: 
// Module Name: invShiftRows_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module invShiftRows_tb;

reg [127:0] in;
wire [127:0] out;	


invShiftRows m (in,out);

initial begin
	$monitor("input= %H , output= %h",in,out);
    in = 128'hd42711ae_e0bf98f1_b8b45de5_1e415230;
    #10;
	//in = 128'h_7ad5fda789ef4e272bca100b3d9ff59f;
    //#10;
    $finish;
end
endmodule
