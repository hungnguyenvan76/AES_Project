`timescale 1ns / 1ps

module invShiftRows_tb;

reg [127:0] in;
wire [127:0] out;	


invShiftRows m (in,out);

initial begin
	$monitor("input= %H , output= %h",in,out);
    in = 128'hd4bf5d30_e0b452ae_b84111f1_1e2798e5;
    #10;
	//in = 128'h_7ad5fda789ef4e272bca100b3d9ff59f;
    //#10;
    $finish;
end
endmodule
